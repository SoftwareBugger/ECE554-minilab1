module Multiplication
#()
(
    input [7:0] 
)